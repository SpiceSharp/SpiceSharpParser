﻿Test
I1 1 0 AC 1
R1 1 0 10
.TRAN 0.1 1.5
.AC LIN 1000 1 1000
.END