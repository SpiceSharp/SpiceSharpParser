﻿Lossless transmission line parse test circuit
T1 1 2 3 4 z0 = 230 Td = 120ns
T2 1 2 3 4 z0=250 f=2.6MEG
T3 1 2 3 4 z0=250 f=2.6MEG m = 10
.END
