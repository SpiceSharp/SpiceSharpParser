﻿ArbitraryBehavioral source
B1 1 0 v = {10 * 10}
R1 1 0 10
.SAVE V(1,0)
.OP
.END